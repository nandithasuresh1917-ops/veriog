module fa 
endmodule
