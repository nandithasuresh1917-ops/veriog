module fa 
